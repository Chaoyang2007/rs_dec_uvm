
`define D #0.2//ns // unblocking delay
`define WIDTH 64 // data with
`define N 198 // size of FEC block
`define K 194 // size of data + syncbit
`define T 2   // error correction ability
`define M 12  // number of symbols in a block, 128b(16B) per symbol
`define PERIOD 2

`define UNBLOCKING_DELAY #0.2 // ns, unblocking delay
`define DATA_WIDTH 64 // data width
`define FEC_BLOCK_SIZE 198 // size of FEC block
`define DATA_SYNC_SIZE 194 // size of data + sync bit
`define ERROR_CORRECTION_ABILITY 2 // error correction ability
`define SYMBOLS_IN_BLOCK 12 // number of symbols in a block, 128b (16B) per symbol
`define CLOCK_PERIOD 2 // clock period
